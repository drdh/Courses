`timescale 1 ns / 1 ps

module liangzhu_player (
	clk,
	i_button_n,
	o_audio
);

input clk;
input i_button_n;
output o_audio;

reg [23:0] counter_4Hz;
reg [23:0] counter_6MHz;
reg [13:0] count;
reg [13:0] origin;
reg audio_reg;
reg clk_6MHz;
reg clk_4Hz;
reg [4:0] note;
reg [10:0] len;

assign o_audio = i_button_n ?  1'b1 : audio_reg;

always @ (posedge clk) begin
	counter_6MHz <= counter_6MHz + 1'b1;
	if (counter_6MHz == 1) begin
		clk_6MHz = ~clk_6MHz;
		counter_6MHz <= 24'b0;
	end
end

always @ (posedge clk) begin
	counter_4Hz <= counter_4Hz + 1'b1;
	if (counter_4Hz == 2999999) begin	
		clk_4Hz = ~clk_4Hz;
		counter_4Hz <= 24'b0;
	end
end

always @ (posedge clk_6MHz) begin
    if(count == 16383) begin
        count = origin;
        audio_reg = ~audio_reg;
    end else
		count = count + 1;
end


always @ (posedge clk_4Hz) begin
	case (note)
		'd0: origin <= 'd16383;h
		'd1: origin <= 'd4916;
		'd2: origin <= 'd6168;
		'd3: origin <= 'd7281;
		'd4: origin <= 'd7791;
		'd5: origin <= 'd8730;
		'd6: origin <= 'd9565;
		'd7: origin <= 'd10310;
		'd8: origin <= 'd010647;
		'd9: origin <= 'd011272;
		'd10: origin <= 'd011831;
		'd11: origin <= 'd012087;
		'd12: origin <= 'd012556;
		'd13: origin <= 'd012974;
		'd14: origin <= 'd013346;
		'd15: origin <= 'd13516;
		'd16: origin <= 'd13829;
		'd17: origin <= 'd14108;
		'd18: origin <= 'd11535;
		'd19: origin <= 'd14470;
		'd20: origin <= 'd14678;
		'd21: origin <= 'd14864;
		default: origin <= 'd011111;
    endcase             
end

always @ (posedge clk_4Hz) begin
	if (len == 958)
		len <= 0;
    else
		len <= len + 1;
	case (len)
		0 :note <= 0;
1 :note <= 0;
2 :note <= 0;
3 :note <= 0;
4 :note <= 0;
5 :note <= 0;
6 :note <= 0;
7 :note <= 0;
8 :note <= 0;
9 :note <= 0;
10 :note <= 0;
11 :note <= 0;
12 :note <= 8;
13 :note <= 8;
14 :note <= 7;
15 :note <= 7;
16 :note <= 6;
17 :note <= 6;
18 :note <= 6;
19 :note <= 6;
20 :note <= 10;
21 :note <= 10;
22 :note <= 10;
23 :note <= 10;
24 :note <= 10;
25 :note <= 10;
26 :note <= 10;
27 :note <= 10;
28 :note <= 8;
29 :note <= 8;
30 :note <= 6;
31 :note <= 6;
32 :note <= 7;
33 :note <= 7;
34 :note <= 7;
35 :note <= 7;
36 :note <= 11;
37 :note <= 11;
38 :note <= 11;
39 :note <= 11;
40 :note <= 10;
41 :note <= 10;
42 :note <= 9;
43 :note <= 9;
44 :note <= 9;
45 :note <= 9;
46 :note <= 9;
47 :note <= 9;
48 :note <= 8;
49 :note <= 8;
50 :note <= 9;
51 :note <= 9;
52 :note <= 8;
53 :note <= 8;
54 :note <= 9;
55 :note <= 9;
56 :note <= 10;
57 :note <= 10;
58 :note <= 10;
59 :note <= 10;
60 :note <= 8;
61 :note <= 8;
62 :note <= 7;
63 :note <= 7;
64 :note <= 6;
65 :note <= 6;
66 :note <= 6;
67 :note <= 6;
68 :note <= 9;
69 :note <= 9;
70 :note <= 9;
71 :note <= 9;
72 :note <= 8;
73 :note <= 8;
74 :note <= 7;
75 :note <= 7;
76 :note <= 0;
77 :note <= 0;
78 :note <= 6;
79 :note <= 7;
80 :note <= 8;
81 :note <= 8;
82 :note <= 8;
83 :note <= 8;
84 :note <= 6;
85 :note <= 6;
86 :note <= 6;
87 :note <= 6;
88 :note <= 10;
89 :note <= 10;
90 :note <= 10;
91 :note <= 10;
92 :note <= 8;
93 :note <= 8;
94 :note <= 8;
95 :note <= 8;
96 :note <= 9;
97 :note <= 9;
98 :note <= 9;
99 :note <= 9;
100 :note <= 13;
101 :note <= 13;
102 :note <= 13;
103 :note <= 13;
104 :note <= 12;
105 :note <= 12;
106 :note <= 12;
107 :note <= 12;
108 :note <= 11;
109 :note <= 11;
110 :note <= 10;
111 :note <= 9;
112 :note <= 10;
113 :note <= 10;
114 :note <= 10;
115 :note <= 10;
116 :note <= 10;
117 :note <= 10;
118 :note <= 10;
119 :note <= 10;
120 :note <= 10;
121 :note <= 10;
122 :note <= 10;
123 :note <= 10;
124 :note <= 10;
125 :note <= 10;
126 :note <= 10;
127 :note <= 10;
128 :note <= 10;
129 :note <= 10;
130 :note <= 10;
131 :note <= 10;
132 :note <= 10;
133 :note <= 10;
134 :note <= 10;
135 :note <= 10;
136 :note <= 0;
137 :note <= 0;
138 :note <= 0;
139 :note <= 0;
140 :note <= 8;
141 :note <= 8;
142 :note <= 7;
143 :note <= 7;
144 :note <= 6;
145 :note <= 6;
146 :note <= 6;
147 :note <= 6;
148 :note <= 10;
149 :note <= 10;
150 :note <= 10;
151 :note <= 10;
152 :note <= 10;
153 :note <= 10;
154 :note <= 10;
155 :note <= 10;
156 :note <= 8;
157 :note <= 8;
158 :note <= 6;
159 :note <= 6;
160 :note <= 7;
161 :note <= 7;
162 :note <= 7;
163 :note <= 7;
164 :note <= 11;
165 :note <= 11;
166 :note <= 11;
167 :note <= 11;
168 :note <= 10;
169 :note <= 10;
170 :note <= 9;
171 :note <= 9;
172 :note <= 9;
173 :note <= 9;
174 :note <= 9;
175 :note <= 9;
176 :note <= 8;
177 :note <= 8;
178 :note <= 9;
179 :note <= 9;
180 :note <= 8;
181 :note <= 8;
182 :note <= 9;
183 :note <= 9;
184 :note <= 10;
185 :note <= 10;
186 :note <= 10;
187 :note <= 10;
188 :note <= 8;
189 :note <= 8;
190 :note <= 7;
191 :note <= 7;
192 :note <= 6;
193 :note <= 6;
194 :note <= 6;
195 :note <= 6;
196 :note <= 9;
197 :note <= 9;
198 :note <= 9;
199 :note <= 9;
200 :note <= 8;
201 :note <= 8;
202 :note <= 7;
203 :note <= 7;
204 :note <= 0;
205 :note <= 0;
206 :note <= 6;
207 :note <= 7;
208 :note <= 8;
209 :note <= 8;
210 :note <= 8;
211 :note <= 8;
212 :note <= 6;
213 :note <= 6;
214 :note <= 6;
215 :note <= 6;
216 :note <= 10;
217 :note <= 10;
218 :note <= 10;
219 :note <= 10;
220 :note <= 8;
221 :note <= 8;
222 :note <= 8;
223 :note <= 8;
224 :note <= 9;
225 :note <= 9;
226 :note <= 9;
227 :note <= 9;
228 :note <= 13;
229 :note <= 13;
230 :note <= 13;
231 :note <= 13;
232 :note <= 12;
233 :note <= 12;
234 :note <= 12;
235 :note <= 12;
236 :note <= 11;
237 :note <= 11;
238 :note <= 10;
239 :note <= 9;
240 :note <= 10;
241 :note <= 10;
242 :note <= 10;
243 :note <= 10;
244 :note <= 10;
245 :note <= 10;
246 :note <= 10;
247 :note <= 10;
248 :note <= 10;
249 :note <= 10;
250 :note <= 10;
251 :note <= 10;
252 :note <= 10;
253 :note <= 10;
254 :note <= 10;
255 :note <= 10;
256 :note <= 10;
257 :note <= 10;
258 :note <= 10;
259 :note <= 10;
260 :note <= 10;
261 :note <= 10;
262 :note <= 10;
263 :note <= 10;
264 :note <= 0;
265 :note <= 0;
266 :note <= 0;
267 :note <= 0;
268 :note <= 10;
269 :note <= 10;
270 :note <= 10;
271 :note <= 10;
272 :note <= 15;
273 :note <= 15;
274 :note <= 15;
275 :note <= 15;
276 :note <= 13;
277 :note <= 13;
278 :note <= 13;
279 :note <= 13;
280 :note <= 13;
281 :note <= 13;
282 :note <= 12;
283 :note <= 12;
284 :note <= 13;
285 :note <= 13;
286 :note <= 15;
287 :note <= 15;
288 :note <= 14;
289 :note <= 14;
290 :note <= 13;
291 :note <= 13;
292 :note <= 13;
293 :note <= 13;
294 :note <= 12;
295 :note <= 12;
296 :note <= 12;
297 :note <= 12;
298 :note <= 12;
299 :note <= 12;
300 :note <= 12;
301 :note <= 12;
302 :note <= 12;
303 :note <= 12;
304 :note <= 13;
305 :note <= 13;
306 :note <= 13;
307 :note <= 13;
308 :note <= 8;
309 :note <= 8;
310 :note <= 9;
311 :note <= 9;
312 :note <= 9;
313 :note <= 9;
314 :note <= 8;
315 :note <= 8;
316 :note <= 9;
317 :note <= 9;
318 :note <= 10;
319 :note <= 10;
320 :note <= 10;
321 :note <= 10;
322 :note <= 10;
323 :note <= 10;
324 :note <= 10;
325 :note <= 10;
326 :note <= 10;
327 :note <= 0;
328 :note <= 0;
329 :note <= 8;
330 :note <= 8;
331 :note <= 9;
332 :note <= 9;
333 :note <= 10;
334 :note <= 10;
335 :note <= 11;
336 :note <= 11;
337 :note <= 11;
338 :note <= 11;
339 :note <= 10;
340 :note <= 10;
341 :note <= 9;
342 :note <= 9;
343 :note <= 9;
344 :note <= 9;
345 :note <= 9;
346 :note <= 9;
347 :note <= 9;
348 :note <= 9;
349 :note <= 9;
350 :note <= 9;
351 :note <= 13;
352 :note <= 13;
353 :note <= 13;
354 :note <= 13;
355 :note <= 12;
356 :note <= 12;
357 :note <= 11;
358 :note <= 11;
359 :note <= 12;
360 :note <= 12;
361 :note <= 13;
362 :note <= 13;
363 :note <= 13;
364 :note <= 13;
365 :note <= 14;
366 :note <= 14;
367 :note <= 14;
368 :note <= 14;
369 :note <= 14;
370 :note <= 14;
371 :note <= 14;
372 :note <= 14;
373 :note <= 14;
374 :note <= 14;
375 :note <= 14;
376 :note <= 14;
377 :note <= 14;
378 :note <= 14;
379 :note <= 14;
380 :note <= 14;
381 :note <= 14;
382 :note <= 14;
383 :note <= 14;
384 :note <= 14;
385 :note <= 14;
386 :note <= 14;
387 :note <= 14;
388 :note <= 14;
389 :note <= 14;
390 :note <= 14;
391 :note <= 0;
392 :note <= 0;
393 :note <= 0;
394 :note <= 0;
395 :note <= 8;
396 :note <= 8;
397 :note <= 7;
398 :note <= 7;
399 :note <= 6;
400 :note <= 6;
401 :note <= 6;
402 :note <= 6;
403 :note <= 10;
404 :note <= 10;
405 :note <= 10;
406 :note <= 10;
407 :note <= 10;
408 :note <= 10;
409 :note <= 10;
410 :note <= 10;
411 :note <= 8;
412 :note <= 8;
413 :note <= 6;
414 :note <= 6;
415 :note <= 7;
416 :note <= 7;
417 :note <= 7;
418 :note <= 7;
419 :note <= 11;
420 :note <= 11;
421 :note <= 11;
422 :note <= 11;
423 :note <= 10;
424 :note <= 10;
425 :note <= 9;
426 :note <= 9;
427 :note <= 9;
428 :note <= 9;
429 :note <= 9;
430 :note <= 9;
431 :note <= 8;
432 :note <= 8;
433 :note <= 9;
434 :note <= 9;
435 :note <= 8;
436 :note <= 8;
437 :note <= 9;
438 :note <= 9;
439 :note <= 10;
440 :note <= 10;
441 :note <= 10;
442 :note <= 10;
443 :note <= 11;
444 :note <= 11;
445 :note <= 12;
446 :note <= 12;
447 :note <= 13;
448 :note <= 13;
449 :note <= 13;
450 :note <= 13;
451 :note <= 15;
452 :note <= 15;
453 :note <= 15;
454 :note <= 15;
455 :note <= 14;
456 :note <= 14;
457 :note <= 12;
458 :note <= 12;
459 :note <= 12;
460 :note <= 12;
461 :note <= 13;
462 :note <= 13;
463 :note <= 13;
464 :note <= 13;
465 :note <= 13;
466 :note <= 13;
467 :note <= 13;
468 :note <= 13;
469 :note <= 13;
470 :note <= 13;
471 :note <= 13;
472 :note <= 13;
473 :note <= 13;
474 :note <= 13;
475 :note <= 13;
476 :note <= 13;
477 :note <= 13;
478 :note <= 13;
479 :note <= 13;
480 :note <= 13;
481 :note <= 13;
482 :note <= 13;
483 :note <= 13;
484 :note <= 13;
485 :note <= 13;
486 :note <= 13;
487 :note <= 0;
488 :note <= 0;
489 :note <= 8;
490 :note <= 8;
491 :note <= 9;
492 :note <= 9;
493 :note <= 10;
494 :note <= 10;
495 :note <= 10;
496 :note <= 10;
497 :note <= 10;
498 :note <= 10;
499 :note <= 10;
500 :note <= 10;
501 :note <= 10;
502 :note <= 10;
503 :note <= 0;
504 :note <= 0;
505 :note <= 4;
506 :note <= 4;
507 :note <= 5;
508 :note <= 5;
509 :note <= 6;
510 :note <= 6;
511 :note <= 6;
512 :note <= 6;
513 :note <= 7;
514 :note <= 7;
515 :note <= 8;
516 :note <= 8;
517 :note <= 9;
518 :note <= 9;
519 :note <= 9;
520 :note <= 9;
521 :note <= 7;
522 :note <= 7;
523 :note <= 7;
524 :note <= 7;
525 :note <= 7;
526 :note <= 7;
527 :note <= 0;
528 :note <= 0;
529 :note <= 0;
530 :note <= 0;
531 :note <= 0;
532 :note <= 0;
533 :note <= 0;
534 :note <= 0;
535 :note <= 0;
536 :note <= 0;
537 :note <= 6;
538 :note <= 6;
539 :note <= 7;
540 :note <= 7;
541 :note <= 8;
542 :note <= 8;
543 :note <= 8;
544 :note <= 8;
545 :note <= 8;
546 :note <= 8;
547 :note <= 8;
548 :note <= 8;
549 :note <= 8;
550 :note <= 8;
551 :note <= 0;
552 :note <= 0;
553 :note <= 8;
554 :note <= 8;
555 :note <= 9;
556 :note <= 9;
557 :note <= 10;
558 :note <= 10;
559 :note <= 10;
560 :note <= 10;
561 :note <= 10;
562 :note <= 10;
563 :note <= 10;
564 :note <= 10;
565 :note <= 10;
566 :note <= 10;
567 :note <= 0;
568 :note <= 0;
569 :note <= 9;
570 :note <= 9;
571 :note <= 10;
572 :note <= 10;
573 :note <= 11;
574 :note <= 12;
575 :note <= 12;
576 :note <= 12;
577 :note <= 12;
578 :note <= 12;
579 :note <= 11;
580 :note <= 11;
581 :note <= 10;
582 :note <= 10;
583 :note <= 10;
584 :note <= 10;
585 :note <= 10;
586 :note <= 10;
587 :note <= 8;
588 :note <= 8;
589 :note <= 7;
590 :note <= 7;
591 :note <= 0;
592 :note <= 0;
593 :note <= 0;
594 :note <= 0;
595 :note <= 0;
596 :note <= 0;
597 :note <= 0;
598 :note <= 0;
599 :note <= 0;
600 :note <= 0;
601 :note <= 0;
602 :note <= 0;
603 :note <= 10;
604 :note <= 10;
605 :note <= 10;
606 :note <= 10;
607 :note <= 15;
608 :note <= 15;
609 :note <= 15;
610 :note <= 15;
611 :note <= 13;
612 :note <= 13;
613 :note <= 13;
614 :note <= 13;
615 :note <= 13;
616 :note <= 13;
617 :note <= 12;
618 :note <= 12;
619 :note <= 13;
620 :note <= 13;
621 :note <= 15;
622 :note <= 15;
623 :note <= 14;
624 :note <= 14;
625 :note <= 13;
626 :note <= 13;
627 :note <= 13;
628 :note <= 13;
629 :note <= 12;
630 :note <= 12;
631 :note <= 12;
632 :note <= 12;
633 :note <= 12;
634 :note <= 12;
635 :note <= 12;
636 :note <= 12;
637 :note <= 12;
638 :note <= 12;
639 :note <= 13;
640 :note <= 13;
641 :note <= 13;
642 :note <= 13;
643 :note <= 8;
644 :note <= 8;
645 :note <= 9;
646 :note <= 9;
647 :note <= 9;
648 :note <= 9;
649 :note <= 8;
650 :note <= 8;
651 :note <= 9;
652 :note <= 9;
653 :note <= 10;
654 :note <= 10;
655 :note <= 10;
656 :note <= 10;
657 :note <= 10;
658 :note <= 10;
659 :note <= 10;
660 :note <= 10;
661 :note <= 10;
662 :note <= 10;
663 :note <= 0;
664 :note <= 0;
665 :note <= 8;
666 :note <= 8;
667 :note <= 9;
668 :note <= 9;
669 :note <= 10;
670 :note <= 10;
671 :note <= 11;
672 :note <= 11;
673 :note <= 11;
674 :note <= 11;
675 :note <= 10;
676 :note <= 10;
677 :note <= 9;
678 :note <= 9;
679 :note <= 9;
680 :note <= 9;
681 :note <= 9;
682 :note <= 9;
683 :note <= 9;
684 :note <= 9;
685 :note <= 9;
686 :note <= 9;
687 :note <= 13;
688 :note <= 13;
689 :note <= 13;
690 :note <= 13;
691 :note <= 12;
692 :note <= 12;
693 :note <= 11;
694 :note <= 11;
695 :note <= 12;
696 :note <= 12;
697 :note <= 13;
698 :note <= 13;
699 :note <= 13;
700 :note <= 13;
701 :note <= 14;
702 :note <= 14;
703 :note <= 14;
704 :note <= 14;
705 :note <= 14;
706 :note <= 14;
707 :note <= 14;
708 :note <= 14;
709 :note <= 14;
710 :note <= 14;
711 :note <= 14;
712 :note <= 14;
713 :note <= 14;
714 :note <= 14;
715 :note <= 14;
716 :note <= 14;
717 :note <= 14;
718 :note <= 14;
719 :note <= 14;
720 :note <= 14;
721 :note <= 14;
722 :note <= 14;
723 :note <= 14;
724 :note <= 14;
725 :note <= 14;
726 :note <= 14;
727 :note <= 0;
728 :note <= 0;
729 :note <= 0;
730 :note <= 0;
731 :note <= 8;
732 :note <= 8;
733 :note <= 7;
734 :note <= 7;
735 :note <= 6;
736 :note <= 6;
737 :note <= 6;
738 :note <= 6;
739 :note <= 10;
740 :note <= 10;
741 :note <= 10;
742 :note <= 10;
743 :note <= 10;
744 :note <= 10;
745 :note <= 10;
746 :note <= 10;
747 :note <= 8;
748 :note <= 8;
749 :note <= 6;
750 :note <= 6;
751 :note <= 7;
752 :note <= 7;
753 :note <= 7;
754 :note <= 7;
755 :note <= 11;
756 :note <= 11;
757 :note <= 11;
758 :note <= 11;
759 :note <= 10;
760 :note <= 10;
761 :note <= 9;
762 :note <= 9;
763 :note <= 9;
764 :note <= 9;
765 :note <= 9;
766 :note <= 9;
767 :note <= 8;
768 :note <= 8;
769 :note <= 9;
770 :note <= 9;
771 :note <= 8;
772 :note <= 8;
773 :note <= 9;
774 :note <= 9;
775 :note <= 10;
776 :note <= 10;
777 :note <= 10;
778 :note <= 10;
779 :note <= 11;
780 :note <= 11;
781 :note <= 12;
782 :note <= 12;
783 :note <= 13;
784 :note <= 13;
785 :note <= 13;
786 :note <= 13;
787 :note <= 15;
788 :note <= 15;
789 :note <= 15;
790 :note <= 15;
791 :note <= 14;
792 :note <= 14;
793 :note <= 12;
794 :note <= 12;
795 :note <= 12;
796 :note <= 12;
797 :note <= 13;
798 :note <= 13;
799 :note <= 13;
800 :note <= 13;
801 :note <= 13;
802 :note <= 13;
803 :note <= 13;
804 :note <= 13;
805 :note <= 13;
806 :note <= 13;
807 :note <= 13;
808 :note <= 13;
809 :note <= 13;
810 :note <= 13;
811 :note <= 13;
812 :note <= 13;
813 :note <= 13;
814 :note <= 13;
815 :note <= 13;
816 :note <= 13;
817 :note <= 13;
818 :note <= 13;
819 :note <= 13;
820 :note <= 13;
821 :note <= 13;
822 :note <= 13;
823 :note <= 13;
824 :note <= 13;
825 :note <= 13;
826 :note <= 13;
827 :note <= 13;
828 :note <= 13;
829 :note <= 13;
830 :note <= 13;
831 :note <= 13;
832 :note <= 13;
833 :note <= 13;
834 :note <= 13;
835 :note <= 13;
836 :note <= 13;
837 :note <= 13;
838 :note <= 13;
839 :note <= 13;
840 :note <= 13;
841 :note <= 13;
842 :note <= 13;
843 :note <= 13;
844 :note <= 13;
845 :note <= 13;
846 :note <= 13;
847 :note <= 12;
848 :note <= 12;
849 :note <= 12;
850 :note <= 12;
851 :note <= 12;
852 :note <= 12;
853 :note <= 11;
854 :note <= 11;
855 :note <= 11;
856 :note <= 11;
857 :note <= 10;
858 :note <= 10;
859 :note <= 9;
860 :note <= 9;
861 :note <= 10;
862 :note <= 10;
863 :note <= 10;
864 :note <= 10;
865 :note <= 10;
866 :note <= 10;
867 :note <= 10;
868 :note <= 10;
869 :note <= 10;
870 :note <= 10;
871 :note <= 10;
872 :note <= 10;
873 :note <= 10;
874 :note <= 10;
875 :note <= 10;
876 :note <= 10;
877 :note <= 10;
878 :note <= 10;
879 :note <= 10;
880 :note <= 10;
881 :note <= 10;
882 :note <= 10;
883 :note <= 10;
884 :note <= 10;
885 :note <= 10;
886 :note <= 10;
887 :note <= 0;
888 :note <= 0;
889 :note <= 11;
890 :note <= 11;
891 :note <= 12;
892 :note <= 12;
893 :note <= 13;
894 :note <= 13;
895 :note <= 13;
896 :note <= 13;
897 :note <= 13;
898 :note <= 13;
899 :note <= 13;
900 :note <= 13;
901 :note <= 13;
902 :note <= 13;
903 :note <= 13;
904 :note <= 13;
905 :note <= 13;
906 :note <= 13;
907 :note <= 13;
908 :note <= 13;
909 :note <= 13;
910 :note <= 13;
911 :note <= 0;
912 :note <= 0;
913 :note <= 0;
914 :note <= 0;
915 :note <= 0;
916 :note <= 0;
917 :note <= 0;
918 :note <= 0;
919 :note <= 0;
920 :note <= 0;
921 :note <= 0;
922 :note <= 0;
923 :note <= 0;
924 :note <= 0;
925 :note <= 0;
926 :note <= 0;
927 :note <= 0;
928 :note <= 0;
929 :note <= 0;
930 :note <= 0;
931 :note <= 0;
932 :note <= 0;
933 :note <= 0;
934 :note <= 0;
935 :note <= 0;
936 :note <= 0;
937 :note <= 0;
938 :note <= 0;
939 :note <= 0;
940 :note <= 0;
941 :note <= 12;
942 :note <= 12;
943 :note <= 13;
944 :note <= 13;
945 :note <= 10;
946 :note <= 10;
947 :note <= 11;
948 :note <= 11;
949 :note <= 9;
950 :note <= 9;
951 :note <= 10;
952 :note <= 10;
953 :note <= 7;
954 :note <= 7;
955 :note <= 8;
956 :note <= 8;
957 :note <= 6;
958 :note <= 6;

	endcase            
end
endmodule