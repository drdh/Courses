
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg  [31:0] ram_cell[0:768-1];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h80f98528;
    ram_cell[       1] = 32'h0;  // 32'hb5aa38c7;
    ram_cell[       2] = 32'h0;  // 32'h0a781dcf;
    ram_cell[       3] = 32'h0;  // 32'h8ff1298f;
    ram_cell[       4] = 32'h0;  // 32'he2aaa08b;
    ram_cell[       5] = 32'h0;  // 32'h2a5828ad;
    ram_cell[       6] = 32'h0;  // 32'h090831c1;
    ram_cell[       7] = 32'h0;  // 32'h966b30cd;
    ram_cell[       8] = 32'h0;  // 32'h40770150;
    ram_cell[       9] = 32'h0;  // 32'h1f0515a7;
    ram_cell[      10] = 32'h0;  // 32'h3654c9ae;
    ram_cell[      11] = 32'h0;  // 32'h192b5670;
    ram_cell[      12] = 32'h0;  // 32'h02f71f5a;
    ram_cell[      13] = 32'h0;  // 32'h52adf15f;
    ram_cell[      14] = 32'h0;  // 32'h3f783f27;
    ram_cell[      15] = 32'h0;  // 32'ha908f4ea;
    ram_cell[      16] = 32'h0;  // 32'he9c33f7b;
    ram_cell[      17] = 32'h0;  // 32'h26dcf3d6;
    ram_cell[      18] = 32'h0;  // 32'hab815621;
    ram_cell[      19] = 32'h0;  // 32'h996186ab;
    ram_cell[      20] = 32'h0;  // 32'h1d93354c;
    ram_cell[      21] = 32'h0;  // 32'h6e54e8fd;
    ram_cell[      22] = 32'h0;  // 32'hf9a7a9e2;
    ram_cell[      23] = 32'h0;  // 32'h7daec384;
    ram_cell[      24] = 32'h0;  // 32'hc6c94b44;
    ram_cell[      25] = 32'h0;  // 32'h722077b2;
    ram_cell[      26] = 32'h0;  // 32'h5b6c3ad6;
    ram_cell[      27] = 32'h0;  // 32'h6c02e112;
    ram_cell[      28] = 32'h0;  // 32'h8aa4002c;
    ram_cell[      29] = 32'h0;  // 32'h6e046c58;
    ram_cell[      30] = 32'h0;  // 32'h01923057;
    ram_cell[      31] = 32'h0;  // 32'hec8fbece;
    ram_cell[      32] = 32'h0;  // 32'h3b2b1057;
    ram_cell[      33] = 32'h0;  // 32'h9ef3d295;
    ram_cell[      34] = 32'h0;  // 32'haacefc60;
    ram_cell[      35] = 32'h0;  // 32'ha3293c25;
    ram_cell[      36] = 32'h0;  // 32'h32b7effa;
    ram_cell[      37] = 32'h0;  // 32'h980dfe9d;
    ram_cell[      38] = 32'h0;  // 32'hdc7a6ccc;
    ram_cell[      39] = 32'h0;  // 32'h6ba4f1fe;
    ram_cell[      40] = 32'h0;  // 32'h0a8cbc9b;
    ram_cell[      41] = 32'h0;  // 32'h849a5ff8;
    ram_cell[      42] = 32'h0;  // 32'h797412a1;
    ram_cell[      43] = 32'h0;  // 32'hfdee6c5d;
    ram_cell[      44] = 32'h0;  // 32'h6172515d;
    ram_cell[      45] = 32'h0;  // 32'hacf2c361;
    ram_cell[      46] = 32'h0;  // 32'hf5bad54c;
    ram_cell[      47] = 32'h0;  // 32'hda1158d6;
    ram_cell[      48] = 32'h0;  // 32'h6037a801;
    ram_cell[      49] = 32'h0;  // 32'h67cbc248;
    ram_cell[      50] = 32'h0;  // 32'h1fbb72ce;
    ram_cell[      51] = 32'h0;  // 32'he0154852;
    ram_cell[      52] = 32'h0;  // 32'hec89bb8e;
    ram_cell[      53] = 32'h0;  // 32'h09f4537e;
    ram_cell[      54] = 32'h0;  // 32'h36308eca;
    ram_cell[      55] = 32'h0;  // 32'he6d034d8;
    ram_cell[      56] = 32'h0;  // 32'haa32e931;
    ram_cell[      57] = 32'h0;  // 32'h25688439;
    ram_cell[      58] = 32'h0;  // 32'h4897f2d6;
    ram_cell[      59] = 32'h0;  // 32'h66f24a08;
    ram_cell[      60] = 32'h0;  // 32'h37328bba;
    ram_cell[      61] = 32'h0;  // 32'h1e3aac4d;
    ram_cell[      62] = 32'h0;  // 32'haea5d0fa;
    ram_cell[      63] = 32'h0;  // 32'hb4145207;
    ram_cell[      64] = 32'h0;  // 32'h3bd8c9c9;
    ram_cell[      65] = 32'h0;  // 32'he8d039e2;
    ram_cell[      66] = 32'h0;  // 32'hae185645;
    ram_cell[      67] = 32'h0;  // 32'h9fcd3b69;
    ram_cell[      68] = 32'h0;  // 32'h8dd3b876;
    ram_cell[      69] = 32'h0;  // 32'h18cf2b47;
    ram_cell[      70] = 32'h0;  // 32'h47ab80a0;
    ram_cell[      71] = 32'h0;  // 32'h81d72cae;
    ram_cell[      72] = 32'h0;  // 32'h1dd37956;
    ram_cell[      73] = 32'h0;  // 32'haca539bb;
    ram_cell[      74] = 32'h0;  // 32'h8f73db13;
    ram_cell[      75] = 32'h0;  // 32'h803230f2;
    ram_cell[      76] = 32'h0;  // 32'h01d8dfd1;
    ram_cell[      77] = 32'h0;  // 32'h700063d0;
    ram_cell[      78] = 32'h0;  // 32'hf958f65f;
    ram_cell[      79] = 32'h0;  // 32'h9a2a6e39;
    ram_cell[      80] = 32'h0;  // 32'h5fc42bc2;
    ram_cell[      81] = 32'h0;  // 32'h636898f3;
    ram_cell[      82] = 32'h0;  // 32'hf9dda6ca;
    ram_cell[      83] = 32'h0;  // 32'hfd2491ee;
    ram_cell[      84] = 32'h0;  // 32'h6dad0f46;
    ram_cell[      85] = 32'h0;  // 32'ha5d6b8a9;
    ram_cell[      86] = 32'h0;  // 32'h2104a6a6;
    ram_cell[      87] = 32'h0;  // 32'hedc14bc7;
    ram_cell[      88] = 32'h0;  // 32'hf14cd0c8;
    ram_cell[      89] = 32'h0;  // 32'h5139c818;
    ram_cell[      90] = 32'h0;  // 32'hc137e677;
    ram_cell[      91] = 32'h0;  // 32'hc34fa341;
    ram_cell[      92] = 32'h0;  // 32'h25ca6eec;
    ram_cell[      93] = 32'h0;  // 32'hb25ec42d;
    ram_cell[      94] = 32'h0;  // 32'hbd8782d9;
    ram_cell[      95] = 32'h0;  // 32'haa364d94;
    ram_cell[      96] = 32'h0;  // 32'h343c5048;
    ram_cell[      97] = 32'h0;  // 32'hab0ade70;
    ram_cell[      98] = 32'h0;  // 32'h1e48cbfe;
    ram_cell[      99] = 32'h0;  // 32'h79c9c445;
    ram_cell[     100] = 32'h0;  // 32'h852dc5d4;
    ram_cell[     101] = 32'h0;  // 32'h38354519;
    ram_cell[     102] = 32'h0;  // 32'hbf6512fc;
    ram_cell[     103] = 32'h0;  // 32'h22e3fc6f;
    ram_cell[     104] = 32'h0;  // 32'h580514dd;
    ram_cell[     105] = 32'h0;  // 32'had459305;
    ram_cell[     106] = 32'h0;  // 32'h5bdebe63;
    ram_cell[     107] = 32'h0;  // 32'hf4eb1dd3;
    ram_cell[     108] = 32'h0;  // 32'hcc900747;
    ram_cell[     109] = 32'h0;  // 32'ha757dc70;
    ram_cell[     110] = 32'h0;  // 32'h3e66fa34;
    ram_cell[     111] = 32'h0;  // 32'h4779cf72;
    ram_cell[     112] = 32'h0;  // 32'h56da78f4;
    ram_cell[     113] = 32'h0;  // 32'h5c12191b;
    ram_cell[     114] = 32'h0;  // 32'hf19556d1;
    ram_cell[     115] = 32'h0;  // 32'hc572dab5;
    ram_cell[     116] = 32'h0;  // 32'hf1418517;
    ram_cell[     117] = 32'h0;  // 32'hf1feee8d;
    ram_cell[     118] = 32'h0;  // 32'h5a0ccb13;
    ram_cell[     119] = 32'h0;  // 32'h1556017f;
    ram_cell[     120] = 32'h0;  // 32'h8d67a106;
    ram_cell[     121] = 32'h0;  // 32'h9774c9bc;
    ram_cell[     122] = 32'h0;  // 32'he186d0bf;
    ram_cell[     123] = 32'h0;  // 32'ha4f27b4f;
    ram_cell[     124] = 32'h0;  // 32'h2cccdbb4;
    ram_cell[     125] = 32'h0;  // 32'hbb4ebbe7;
    ram_cell[     126] = 32'h0;  // 32'h94ee994a;
    ram_cell[     127] = 32'h0;  // 32'h29719bd6;
    ram_cell[     128] = 32'h0;  // 32'hd1a57ada;
    ram_cell[     129] = 32'h0;  // 32'h96bde61e;
    ram_cell[     130] = 32'h0;  // 32'h5c8099d6;
    ram_cell[     131] = 32'h0;  // 32'hefaf9a9f;
    ram_cell[     132] = 32'h0;  // 32'hb6a4941e;
    ram_cell[     133] = 32'h0;  // 32'h221d420e;
    ram_cell[     134] = 32'h0;  // 32'h22fb6993;
    ram_cell[     135] = 32'h0;  // 32'h1d90ef70;
    ram_cell[     136] = 32'h0;  // 32'hc84ba9f6;
    ram_cell[     137] = 32'h0;  // 32'h8e0e621a;
    ram_cell[     138] = 32'h0;  // 32'h110468e3;
    ram_cell[     139] = 32'h0;  // 32'h60c6c354;
    ram_cell[     140] = 32'h0;  // 32'h0411b39f;
    ram_cell[     141] = 32'h0;  // 32'h448ade5c;
    ram_cell[     142] = 32'h0;  // 32'h2bca6d9b;
    ram_cell[     143] = 32'h0;  // 32'h15461576;
    ram_cell[     144] = 32'h0;  // 32'h066b0f1d;
    ram_cell[     145] = 32'h0;  // 32'he4a5f481;
    ram_cell[     146] = 32'h0;  // 32'h337ee658;
    ram_cell[     147] = 32'h0;  // 32'h1900d3c3;
    ram_cell[     148] = 32'h0;  // 32'h8f53a25c;
    ram_cell[     149] = 32'h0;  // 32'h8545666c;
    ram_cell[     150] = 32'h0;  // 32'h61d9f55a;
    ram_cell[     151] = 32'h0;  // 32'h6109bbbf;
    ram_cell[     152] = 32'h0;  // 32'hb0c4a297;
    ram_cell[     153] = 32'h0;  // 32'he71a44b9;
    ram_cell[     154] = 32'h0;  // 32'h6cea1e4e;
    ram_cell[     155] = 32'h0;  // 32'hd3f6f704;
    ram_cell[     156] = 32'h0;  // 32'h75787a8c;
    ram_cell[     157] = 32'h0;  // 32'h0d52dacf;
    ram_cell[     158] = 32'h0;  // 32'h5785f584;
    ram_cell[     159] = 32'h0;  // 32'hf3d920c1;
    ram_cell[     160] = 32'h0;  // 32'h2dcd5899;
    ram_cell[     161] = 32'h0;  // 32'h5e6bf2ce;
    ram_cell[     162] = 32'h0;  // 32'hbdb48161;
    ram_cell[     163] = 32'h0;  // 32'h09c3d7cc;
    ram_cell[     164] = 32'h0;  // 32'h9f83de4c;
    ram_cell[     165] = 32'h0;  // 32'h83f9438d;
    ram_cell[     166] = 32'h0;  // 32'ha78fb8a5;
    ram_cell[     167] = 32'h0;  // 32'h50343ebb;
    ram_cell[     168] = 32'h0;  // 32'hd0022d17;
    ram_cell[     169] = 32'h0;  // 32'h5e686aeb;
    ram_cell[     170] = 32'h0;  // 32'h8e941a59;
    ram_cell[     171] = 32'h0;  // 32'h0afacb1c;
    ram_cell[     172] = 32'h0;  // 32'h718c5dbb;
    ram_cell[     173] = 32'h0;  // 32'hcd123a29;
    ram_cell[     174] = 32'h0;  // 32'h09c858d6;
    ram_cell[     175] = 32'h0;  // 32'h1ced3507;
    ram_cell[     176] = 32'h0;  // 32'hd8a5f713;
    ram_cell[     177] = 32'h0;  // 32'ha3fc7607;
    ram_cell[     178] = 32'h0;  // 32'hf3177873;
    ram_cell[     179] = 32'h0;  // 32'h13cbe9f8;
    ram_cell[     180] = 32'h0;  // 32'h01c9c50b;
    ram_cell[     181] = 32'h0;  // 32'he332c9df;
    ram_cell[     182] = 32'h0;  // 32'hf2990269;
    ram_cell[     183] = 32'h0;  // 32'hb12e6a8a;
    ram_cell[     184] = 32'h0;  // 32'hb5c1431c;
    ram_cell[     185] = 32'h0;  // 32'h400536c9;
    ram_cell[     186] = 32'h0;  // 32'h9d5f9213;
    ram_cell[     187] = 32'h0;  // 32'h9cc74e52;
    ram_cell[     188] = 32'h0;  // 32'hfd1b0c09;
    ram_cell[     189] = 32'h0;  // 32'hb1f04d4a;
    ram_cell[     190] = 32'h0;  // 32'hf6b9b21d;
    ram_cell[     191] = 32'h0;  // 32'h64df2a5f;
    ram_cell[     192] = 32'h0;  // 32'hbdd71731;
    ram_cell[     193] = 32'h0;  // 32'h6547fe1c;
    ram_cell[     194] = 32'h0;  // 32'h06c6c479;
    ram_cell[     195] = 32'h0;  // 32'hd8e6c6ec;
    ram_cell[     196] = 32'h0;  // 32'h51b5e1cd;
    ram_cell[     197] = 32'h0;  // 32'h73c63594;
    ram_cell[     198] = 32'h0;  // 32'h526e0b66;
    ram_cell[     199] = 32'h0;  // 32'h4f327e3b;
    ram_cell[     200] = 32'h0;  // 32'h6298d50e;
    ram_cell[     201] = 32'h0;  // 32'h6b8699ae;
    ram_cell[     202] = 32'h0;  // 32'h01d1d23b;
    ram_cell[     203] = 32'h0;  // 32'ha1b9958a;
    ram_cell[     204] = 32'h0;  // 32'hef02cccd;
    ram_cell[     205] = 32'h0;  // 32'h08d9eb5c;
    ram_cell[     206] = 32'h0;  // 32'hed4519ba;
    ram_cell[     207] = 32'h0;  // 32'hc926320a;
    ram_cell[     208] = 32'h0;  // 32'h231535f0;
    ram_cell[     209] = 32'h0;  // 32'h51bc8772;
    ram_cell[     210] = 32'h0;  // 32'h18985870;
    ram_cell[     211] = 32'h0;  // 32'h469b434f;
    ram_cell[     212] = 32'h0;  // 32'ha043264b;
    ram_cell[     213] = 32'h0;  // 32'h517333c9;
    ram_cell[     214] = 32'h0;  // 32'h9937e573;
    ram_cell[     215] = 32'h0;  // 32'h2a60316a;
    ram_cell[     216] = 32'h0;  // 32'h4a45454b;
    ram_cell[     217] = 32'h0;  // 32'h3b97c6e5;
    ram_cell[     218] = 32'h0;  // 32'hb21deb10;
    ram_cell[     219] = 32'h0;  // 32'h08e41bc2;
    ram_cell[     220] = 32'h0;  // 32'h7da2d2f5;
    ram_cell[     221] = 32'h0;  // 32'h86af33ea;
    ram_cell[     222] = 32'h0;  // 32'hf883b424;
    ram_cell[     223] = 32'h0;  // 32'h5a68b236;
    ram_cell[     224] = 32'h0;  // 32'h96ac98d1;
    ram_cell[     225] = 32'h0;  // 32'h5402fa94;
    ram_cell[     226] = 32'h0;  // 32'h0fa31028;
    ram_cell[     227] = 32'h0;  // 32'h23292a35;
    ram_cell[     228] = 32'h0;  // 32'h3eff74e6;
    ram_cell[     229] = 32'h0;  // 32'h92efb58a;
    ram_cell[     230] = 32'h0;  // 32'he50fafa6;
    ram_cell[     231] = 32'h0;  // 32'h0fe95aad;
    ram_cell[     232] = 32'h0;  // 32'haeb8201a;
    ram_cell[     233] = 32'h0;  // 32'hbdef6ce2;
    ram_cell[     234] = 32'h0;  // 32'h13a730a2;
    ram_cell[     235] = 32'h0;  // 32'h5abd1ca3;
    ram_cell[     236] = 32'h0;  // 32'h250330bb;
    ram_cell[     237] = 32'h0;  // 32'hfe9e53dc;
    ram_cell[     238] = 32'h0;  // 32'he858e5b0;
    ram_cell[     239] = 32'h0;  // 32'h3482d88b;
    ram_cell[     240] = 32'h0;  // 32'hc47d1eb6;
    ram_cell[     241] = 32'h0;  // 32'h35916274;
    ram_cell[     242] = 32'h0;  // 32'h671bcf54;
    ram_cell[     243] = 32'h0;  // 32'hfa010e93;
    ram_cell[     244] = 32'h0;  // 32'hc90daf08;
    ram_cell[     245] = 32'h0;  // 32'h6d587967;
    ram_cell[     246] = 32'h0;  // 32'h5d485b44;
    ram_cell[     247] = 32'h0;  // 32'hec0e5d01;
    ram_cell[     248] = 32'h0;  // 32'h10f2d4c2;
    ram_cell[     249] = 32'h0;  // 32'h5a28cf06;
    ram_cell[     250] = 32'h0;  // 32'h01bf4f68;
    ram_cell[     251] = 32'h0;  // 32'hff7eabc9;
    ram_cell[     252] = 32'h0;  // 32'h1a9b2034;
    ram_cell[     253] = 32'h0;  // 32'h13d69dbd;
    ram_cell[     254] = 32'h0;  // 32'h37a5b890;
    ram_cell[     255] = 32'h0;  // 32'hf7ae234a;
    // src matrix A
    ram_cell[     256] = 32'h17ebacdc;
    ram_cell[     257] = 32'h3cdd158c;
    ram_cell[     258] = 32'h38768f02;
    ram_cell[     259] = 32'h9d3a8f90;
    ram_cell[     260] = 32'h8e4e5e73;
    ram_cell[     261] = 32'hf6febcd5;
    ram_cell[     262] = 32'h1850136c;
    ram_cell[     263] = 32'hc53f6478;
    ram_cell[     264] = 32'hc1e56e14;
    ram_cell[     265] = 32'h4b557e17;
    ram_cell[     266] = 32'h0bc3611c;
    ram_cell[     267] = 32'h4c520854;
    ram_cell[     268] = 32'hb11a4f88;
    ram_cell[     269] = 32'he254cb7d;
    ram_cell[     270] = 32'h06c5bfcc;
    ram_cell[     271] = 32'h24985b48;
    ram_cell[     272] = 32'h28fc7104;
    ram_cell[     273] = 32'had53bcb5;
    ram_cell[     274] = 32'h60f9f761;
    ram_cell[     275] = 32'h6b443455;
    ram_cell[     276] = 32'hfe7c7727;
    ram_cell[     277] = 32'h2cfe78fa;
    ram_cell[     278] = 32'h2d86fc6c;
    ram_cell[     279] = 32'hf71f4b2a;
    ram_cell[     280] = 32'h2929ce6d;
    ram_cell[     281] = 32'h803a7727;
    ram_cell[     282] = 32'h78733d4b;
    ram_cell[     283] = 32'hb19432d3;
    ram_cell[     284] = 32'hb686acdf;
    ram_cell[     285] = 32'ha6f1b100;
    ram_cell[     286] = 32'h444bf114;
    ram_cell[     287] = 32'ha52c1806;
    ram_cell[     288] = 32'h4d4afc7b;
    ram_cell[     289] = 32'h2304faac;
    ram_cell[     290] = 32'hccb9762b;
    ram_cell[     291] = 32'h8ec705c4;
    ram_cell[     292] = 32'hd833d34f;
    ram_cell[     293] = 32'h0945fb48;
    ram_cell[     294] = 32'h740f834e;
    ram_cell[     295] = 32'h2f9d264f;
    ram_cell[     296] = 32'h11f9a5a5;
    ram_cell[     297] = 32'hdc1016b5;
    ram_cell[     298] = 32'h1d05e00f;
    ram_cell[     299] = 32'he0722f42;
    ram_cell[     300] = 32'hf9a1769b;
    ram_cell[     301] = 32'h667035db;
    ram_cell[     302] = 32'h530daac9;
    ram_cell[     303] = 32'h0a21e6f2;
    ram_cell[     304] = 32'h2f4f70d4;
    ram_cell[     305] = 32'hba507e3f;
    ram_cell[     306] = 32'h073d2e35;
    ram_cell[     307] = 32'h16d225a0;
    ram_cell[     308] = 32'hfa13a14d;
    ram_cell[     309] = 32'h284aa0c2;
    ram_cell[     310] = 32'hfb765f83;
    ram_cell[     311] = 32'hafebf5d2;
    ram_cell[     312] = 32'hf935bc2b;
    ram_cell[     313] = 32'h39c1e245;
    ram_cell[     314] = 32'h65317e4c;
    ram_cell[     315] = 32'hf2ef8840;
    ram_cell[     316] = 32'h58179b0f;
    ram_cell[     317] = 32'ha159d498;
    ram_cell[     318] = 32'h80538878;
    ram_cell[     319] = 32'h8cba6d70;
    ram_cell[     320] = 32'h8f0dc878;
    ram_cell[     321] = 32'h4b9f07a1;
    ram_cell[     322] = 32'h8fa4e5b3;
    ram_cell[     323] = 32'h3e448e15;
    ram_cell[     324] = 32'hb47f8fc9;
    ram_cell[     325] = 32'h97bd9226;
    ram_cell[     326] = 32'hfce09f1e;
    ram_cell[     327] = 32'h69c4a3e2;
    ram_cell[     328] = 32'hd2693b87;
    ram_cell[     329] = 32'h67d5ce88;
    ram_cell[     330] = 32'hf558de51;
    ram_cell[     331] = 32'h8e187fe2;
    ram_cell[     332] = 32'hd3c20923;
    ram_cell[     333] = 32'hc6a6a1f2;
    ram_cell[     334] = 32'hd1956ec6;
    ram_cell[     335] = 32'h2426fc82;
    ram_cell[     336] = 32'hdc630722;
    ram_cell[     337] = 32'hda91ca01;
    ram_cell[     338] = 32'h5c6b1d23;
    ram_cell[     339] = 32'h38ca64f9;
    ram_cell[     340] = 32'h778c8b42;
    ram_cell[     341] = 32'hcccdbaee;
    ram_cell[     342] = 32'hc40d5fd7;
    ram_cell[     343] = 32'h487c37d9;
    ram_cell[     344] = 32'he59489db;
    ram_cell[     345] = 32'hca20817d;
    ram_cell[     346] = 32'h09c883bd;
    ram_cell[     347] = 32'h11ce6864;
    ram_cell[     348] = 32'hebef4ac4;
    ram_cell[     349] = 32'hfedabac4;
    ram_cell[     350] = 32'hcc034218;
    ram_cell[     351] = 32'hb8f59320;
    ram_cell[     352] = 32'h0a4b3301;
    ram_cell[     353] = 32'h143aa5fa;
    ram_cell[     354] = 32'h142bf273;
    ram_cell[     355] = 32'h8e1d0472;
    ram_cell[     356] = 32'h09346efb;
    ram_cell[     357] = 32'h3e486263;
    ram_cell[     358] = 32'h407d12da;
    ram_cell[     359] = 32'h11b71229;
    ram_cell[     360] = 32'ha03b24d7;
    ram_cell[     361] = 32'hcc0fbdf2;
    ram_cell[     362] = 32'h6fd291a7;
    ram_cell[     363] = 32'h24d054b0;
    ram_cell[     364] = 32'h9e585008;
    ram_cell[     365] = 32'h839600a0;
    ram_cell[     366] = 32'hfc1a7999;
    ram_cell[     367] = 32'h972043f0;
    ram_cell[     368] = 32'h5a20e9fb;
    ram_cell[     369] = 32'h65d31b4e;
    ram_cell[     370] = 32'h938f7ffa;
    ram_cell[     371] = 32'h34931d80;
    ram_cell[     372] = 32'h8d969fea;
    ram_cell[     373] = 32'had72e916;
    ram_cell[     374] = 32'h6fa15486;
    ram_cell[     375] = 32'h435c1120;
    ram_cell[     376] = 32'hf431f1c8;
    ram_cell[     377] = 32'h6eb26634;
    ram_cell[     378] = 32'h0bc4397e;
    ram_cell[     379] = 32'h9f7591f8;
    ram_cell[     380] = 32'hd37f6901;
    ram_cell[     381] = 32'h924fd090;
    ram_cell[     382] = 32'ha00cd77a;
    ram_cell[     383] = 32'hd2b55c75;
    ram_cell[     384] = 32'hdcbca84f;
    ram_cell[     385] = 32'hcf338935;
    ram_cell[     386] = 32'ha4bf57b5;
    ram_cell[     387] = 32'hc833ad0a;
    ram_cell[     388] = 32'h3c8ad560;
    ram_cell[     389] = 32'hd6f81650;
    ram_cell[     390] = 32'h2978b160;
    ram_cell[     391] = 32'h5f2c2a13;
    ram_cell[     392] = 32'h45e46cdb;
    ram_cell[     393] = 32'he9df0311;
    ram_cell[     394] = 32'hc0871b3d;
    ram_cell[     395] = 32'h17905a80;
    ram_cell[     396] = 32'h4a6417f9;
    ram_cell[     397] = 32'hff9039eb;
    ram_cell[     398] = 32'h771ee57c;
    ram_cell[     399] = 32'hb33df806;
    ram_cell[     400] = 32'he7e2ae79;
    ram_cell[     401] = 32'h344a9d3a;
    ram_cell[     402] = 32'h2e77cfa1;
    ram_cell[     403] = 32'h007c292d;
    ram_cell[     404] = 32'hb008e30a;
    ram_cell[     405] = 32'hf96c029f;
    ram_cell[     406] = 32'hf28ed01c;
    ram_cell[     407] = 32'h15f2a958;
    ram_cell[     408] = 32'h5e8ef725;
    ram_cell[     409] = 32'hcff0e3fc;
    ram_cell[     410] = 32'h3e856607;
    ram_cell[     411] = 32'hc15a62d4;
    ram_cell[     412] = 32'hd78f2cf0;
    ram_cell[     413] = 32'h09658252;
    ram_cell[     414] = 32'hadd9b411;
    ram_cell[     415] = 32'hb7f168c2;
    ram_cell[     416] = 32'h093e9ba1;
    ram_cell[     417] = 32'h3a264058;
    ram_cell[     418] = 32'hc2ab1ca8;
    ram_cell[     419] = 32'hcd319d9f;
    ram_cell[     420] = 32'h838c2ca6;
    ram_cell[     421] = 32'hf5ed6c8b;
    ram_cell[     422] = 32'h131bb53d;
    ram_cell[     423] = 32'h548ea1f4;
    ram_cell[     424] = 32'h027e047b;
    ram_cell[     425] = 32'hc39253a7;
    ram_cell[     426] = 32'h59005e5f;
    ram_cell[     427] = 32'h53537099;
    ram_cell[     428] = 32'h531bc454;
    ram_cell[     429] = 32'h1b8ebaa7;
    ram_cell[     430] = 32'hc69c438b;
    ram_cell[     431] = 32'hb3ac1781;
    ram_cell[     432] = 32'hf3a6f6e9;
    ram_cell[     433] = 32'hfcdd5719;
    ram_cell[     434] = 32'h57e774fb;
    ram_cell[     435] = 32'he46ef504;
    ram_cell[     436] = 32'he0c286c1;
    ram_cell[     437] = 32'h149ad19a;
    ram_cell[     438] = 32'h12767ebc;
    ram_cell[     439] = 32'ha06875e6;
    ram_cell[     440] = 32'hd21eb0f0;
    ram_cell[     441] = 32'h38730287;
    ram_cell[     442] = 32'h4bfbf686;
    ram_cell[     443] = 32'habaaf0e8;
    ram_cell[     444] = 32'hab97683b;
    ram_cell[     445] = 32'h7412cef2;
    ram_cell[     446] = 32'h4e9273f0;
    ram_cell[     447] = 32'h405d43e4;
    ram_cell[     448] = 32'h7977ce04;
    ram_cell[     449] = 32'ha84433dd;
    ram_cell[     450] = 32'h4bf1d033;
    ram_cell[     451] = 32'hc3c2632f;
    ram_cell[     452] = 32'hd2aaf394;
    ram_cell[     453] = 32'h781ad9bb;
    ram_cell[     454] = 32'hcf925b65;
    ram_cell[     455] = 32'hf9a732d5;
    ram_cell[     456] = 32'ha94753d4;
    ram_cell[     457] = 32'h0e0a78a0;
    ram_cell[     458] = 32'hd954ffb3;
    ram_cell[     459] = 32'h416922fc;
    ram_cell[     460] = 32'h31caacc7;
    ram_cell[     461] = 32'h2d57761b;
    ram_cell[     462] = 32'hcdfaaf47;
    ram_cell[     463] = 32'h6a634936;
    ram_cell[     464] = 32'hf8bdf63a;
    ram_cell[     465] = 32'hc42c100f;
    ram_cell[     466] = 32'h5cc62a9c;
    ram_cell[     467] = 32'h59916e75;
    ram_cell[     468] = 32'h25353359;
    ram_cell[     469] = 32'h4318cd64;
    ram_cell[     470] = 32'h1c3182bd;
    ram_cell[     471] = 32'hca289743;
    ram_cell[     472] = 32'ha07b4126;
    ram_cell[     473] = 32'hd49b599c;
    ram_cell[     474] = 32'ha43abdcd;
    ram_cell[     475] = 32'hb747125a;
    ram_cell[     476] = 32'h3d6bb293;
    ram_cell[     477] = 32'h112465a0;
    ram_cell[     478] = 32'hfd9eb867;
    ram_cell[     479] = 32'h588dcecd;
    ram_cell[     480] = 32'hfaf10f65;
    ram_cell[     481] = 32'h7010b789;
    ram_cell[     482] = 32'hb6ecbc4f;
    ram_cell[     483] = 32'h5315ebbd;
    ram_cell[     484] = 32'h8713c296;
    ram_cell[     485] = 32'h462b1732;
    ram_cell[     486] = 32'he2d3cbe9;
    ram_cell[     487] = 32'h9d7f78d5;
    ram_cell[     488] = 32'h163c0b55;
    ram_cell[     489] = 32'h041d7052;
    ram_cell[     490] = 32'hc8fe4877;
    ram_cell[     491] = 32'hc7e6858b;
    ram_cell[     492] = 32'h39d8bf91;
    ram_cell[     493] = 32'hc78f8aef;
    ram_cell[     494] = 32'h6b02971e;
    ram_cell[     495] = 32'h0371afcc;
    ram_cell[     496] = 32'h6fbed492;
    ram_cell[     497] = 32'h7294ec14;
    ram_cell[     498] = 32'h33810898;
    ram_cell[     499] = 32'hff398092;
    ram_cell[     500] = 32'h291e73f3;
    ram_cell[     501] = 32'hebef2e20;
    ram_cell[     502] = 32'h7349e823;
    ram_cell[     503] = 32'h65d7ad89;
    ram_cell[     504] = 32'h8c34d607;
    ram_cell[     505] = 32'hc0051a11;
    ram_cell[     506] = 32'h62bdf431;
    ram_cell[     507] = 32'h8ad5fdab;
    ram_cell[     508] = 32'hdc7e8b36;
    ram_cell[     509] = 32'h48d20fd9;
    ram_cell[     510] = 32'h73a85646;
    ram_cell[     511] = 32'h1dd831d0;
    // src matrix B
    ram_cell[     512] = 32'hac5bf5b0;
    ram_cell[     513] = 32'h7ffc5984;
    ram_cell[     514] = 32'h87d401d3;
    ram_cell[     515] = 32'hc235f8f5;
    ram_cell[     516] = 32'hf2e42862;
    ram_cell[     517] = 32'h43fca4e9;
    ram_cell[     518] = 32'h3b725ad8;
    ram_cell[     519] = 32'he2c69e5b;
    ram_cell[     520] = 32'ha2fc877b;
    ram_cell[     521] = 32'hfdf4dd9c;
    ram_cell[     522] = 32'h8e9e66ff;
    ram_cell[     523] = 32'h8f2a3d20;
    ram_cell[     524] = 32'hc1cec1e0;
    ram_cell[     525] = 32'h53670d49;
    ram_cell[     526] = 32'hc821ac03;
    ram_cell[     527] = 32'h31c57613;
    ram_cell[     528] = 32'h1139a1ae;
    ram_cell[     529] = 32'h55894dc7;
    ram_cell[     530] = 32'hc5f9c0cd;
    ram_cell[     531] = 32'hdd94a87d;
    ram_cell[     532] = 32'h70eb0906;
    ram_cell[     533] = 32'h06f5d3b6;
    ram_cell[     534] = 32'h4ec25452;
    ram_cell[     535] = 32'h4e88ecb4;
    ram_cell[     536] = 32'h01d476b2;
    ram_cell[     537] = 32'h4599827e;
    ram_cell[     538] = 32'h07fc65b7;
    ram_cell[     539] = 32'h512bf596;
    ram_cell[     540] = 32'h6eed179a;
    ram_cell[     541] = 32'hb7f5e4d3;
    ram_cell[     542] = 32'hed1bb87c;
    ram_cell[     543] = 32'hc6e576c9;
    ram_cell[     544] = 32'hacbbdcd0;
    ram_cell[     545] = 32'hd341d7e6;
    ram_cell[     546] = 32'h8be2a013;
    ram_cell[     547] = 32'h94afd215;
    ram_cell[     548] = 32'he79013d4;
    ram_cell[     549] = 32'he87b2195;
    ram_cell[     550] = 32'h28686d2c;
    ram_cell[     551] = 32'h37ca951e;
    ram_cell[     552] = 32'h9494eae4;
    ram_cell[     553] = 32'hf675769e;
    ram_cell[     554] = 32'h8f6bc9b0;
    ram_cell[     555] = 32'hd36bb1b6;
    ram_cell[     556] = 32'h067cf203;
    ram_cell[     557] = 32'h7b48ceed;
    ram_cell[     558] = 32'hb05b3451;
    ram_cell[     559] = 32'h1e6613c9;
    ram_cell[     560] = 32'h57b1117a;
    ram_cell[     561] = 32'h8e5949a1;
    ram_cell[     562] = 32'h0280441b;
    ram_cell[     563] = 32'h23814222;
    ram_cell[     564] = 32'h5a4a0039;
    ram_cell[     565] = 32'hefd039ae;
    ram_cell[     566] = 32'h5b2738c1;
    ram_cell[     567] = 32'h7d787d9e;
    ram_cell[     568] = 32'h8e2304d2;
    ram_cell[     569] = 32'hdacf92eb;
    ram_cell[     570] = 32'h13d9e7c5;
    ram_cell[     571] = 32'h0d9aa8b0;
    ram_cell[     572] = 32'hd6df35d0;
    ram_cell[     573] = 32'hcc82c8a7;
    ram_cell[     574] = 32'h5c59fcd5;
    ram_cell[     575] = 32'hdf59da5e;
    ram_cell[     576] = 32'hd8311cfa;
    ram_cell[     577] = 32'h59c73cb6;
    ram_cell[     578] = 32'h0b15ecf5;
    ram_cell[     579] = 32'he1f445be;
    ram_cell[     580] = 32'hd5752527;
    ram_cell[     581] = 32'h04534502;
    ram_cell[     582] = 32'h428ed37e;
    ram_cell[     583] = 32'h77d356f5;
    ram_cell[     584] = 32'h0340764b;
    ram_cell[     585] = 32'he3a77f21;
    ram_cell[     586] = 32'hc5e2f0fe;
    ram_cell[     587] = 32'h12ae3c5f;
    ram_cell[     588] = 32'h9dc635df;
    ram_cell[     589] = 32'ha6071b7d;
    ram_cell[     590] = 32'ha6e3c2b0;
    ram_cell[     591] = 32'hfc9f0d14;
    ram_cell[     592] = 32'h62aa120c;
    ram_cell[     593] = 32'hc9d734c6;
    ram_cell[     594] = 32'hb39efec0;
    ram_cell[     595] = 32'h76554a28;
    ram_cell[     596] = 32'ha6c020b4;
    ram_cell[     597] = 32'hf23fc95e;
    ram_cell[     598] = 32'h30f215fa;
    ram_cell[     599] = 32'h0133e29f;
    ram_cell[     600] = 32'h783b4df6;
    ram_cell[     601] = 32'h39cfef0f;
    ram_cell[     602] = 32'haac5cfd2;
    ram_cell[     603] = 32'hd32efe42;
    ram_cell[     604] = 32'h0be2dd56;
    ram_cell[     605] = 32'hb4c7f652;
    ram_cell[     606] = 32'h0ddd3152;
    ram_cell[     607] = 32'h900b0841;
    ram_cell[     608] = 32'hb5ac4515;
    ram_cell[     609] = 32'h24ebe927;
    ram_cell[     610] = 32'h819a86f5;
    ram_cell[     611] = 32'hb24d4aae;
    ram_cell[     612] = 32'h3f4f4f1b;
    ram_cell[     613] = 32'h7c4b9d4e;
    ram_cell[     614] = 32'hd6148670;
    ram_cell[     615] = 32'h7cc94e77;
    ram_cell[     616] = 32'hb6f90f34;
    ram_cell[     617] = 32'h4bd3a8da;
    ram_cell[     618] = 32'h01da8b3f;
    ram_cell[     619] = 32'hb3b135bd;
    ram_cell[     620] = 32'h4113ddc9;
    ram_cell[     621] = 32'h839b4bdf;
    ram_cell[     622] = 32'hf612e92c;
    ram_cell[     623] = 32'h867a1dc2;
    ram_cell[     624] = 32'hf330ea2b;
    ram_cell[     625] = 32'hc86cfef6;
    ram_cell[     626] = 32'h6a648b28;
    ram_cell[     627] = 32'h159cbb18;
    ram_cell[     628] = 32'he8e1cdea;
    ram_cell[     629] = 32'heb9a7d51;
    ram_cell[     630] = 32'h5a59496b;
    ram_cell[     631] = 32'h64d595f5;
    ram_cell[     632] = 32'hae9196e5;
    ram_cell[     633] = 32'h2fd6337a;
    ram_cell[     634] = 32'hd3a9d58e;
    ram_cell[     635] = 32'h5cabbb56;
    ram_cell[     636] = 32'h5d5bb78c;
    ram_cell[     637] = 32'hd86e995b;
    ram_cell[     638] = 32'hd75fc3e3;
    ram_cell[     639] = 32'h6c3a42dd;
    ram_cell[     640] = 32'h6523934d;
    ram_cell[     641] = 32'h08b2fff0;
    ram_cell[     642] = 32'hcaa0b1ed;
    ram_cell[     643] = 32'hf06cc52f;
    ram_cell[     644] = 32'he7d2392e;
    ram_cell[     645] = 32'hbea4a32c;
    ram_cell[     646] = 32'h09122ee3;
    ram_cell[     647] = 32'h4afde340;
    ram_cell[     648] = 32'h0658dcd8;
    ram_cell[     649] = 32'h6cfe4a4c;
    ram_cell[     650] = 32'h1120ac1f;
    ram_cell[     651] = 32'hf4195a59;
    ram_cell[     652] = 32'ha9b78c7c;
    ram_cell[     653] = 32'h23d9ed93;
    ram_cell[     654] = 32'h7c85ed8e;
    ram_cell[     655] = 32'hbbfaef31;
    ram_cell[     656] = 32'h7725879e;
    ram_cell[     657] = 32'h77055f6e;
    ram_cell[     658] = 32'hfffd6803;
    ram_cell[     659] = 32'hfabb61b0;
    ram_cell[     660] = 32'h8e54b1e8;
    ram_cell[     661] = 32'he454cd3a;
    ram_cell[     662] = 32'h39e94e56;
    ram_cell[     663] = 32'hc76bcbd5;
    ram_cell[     664] = 32'hb5f8ac85;
    ram_cell[     665] = 32'h51957d27;
    ram_cell[     666] = 32'hdebf34d3;
    ram_cell[     667] = 32'hb12fea82;
    ram_cell[     668] = 32'h2b0b745c;
    ram_cell[     669] = 32'hef5a589d;
    ram_cell[     670] = 32'hf7732d3a;
    ram_cell[     671] = 32'h6f569138;
    ram_cell[     672] = 32'h5ed95c31;
    ram_cell[     673] = 32'h0098cff4;
    ram_cell[     674] = 32'h154ca4b8;
    ram_cell[     675] = 32'h7fe759bd;
    ram_cell[     676] = 32'hae227d96;
    ram_cell[     677] = 32'h0c10beed;
    ram_cell[     678] = 32'h2b04d367;
    ram_cell[     679] = 32'h80e8962a;
    ram_cell[     680] = 32'h6e73b562;
    ram_cell[     681] = 32'h7f1fe7a2;
    ram_cell[     682] = 32'h48b46300;
    ram_cell[     683] = 32'h4a819c6f;
    ram_cell[     684] = 32'hceddc7d8;
    ram_cell[     685] = 32'h1bbc0158;
    ram_cell[     686] = 32'h74fffbc6;
    ram_cell[     687] = 32'hbc0d02f8;
    ram_cell[     688] = 32'hfdc6c116;
    ram_cell[     689] = 32'h044dd960;
    ram_cell[     690] = 32'hd4fca643;
    ram_cell[     691] = 32'h29d72cd4;
    ram_cell[     692] = 32'h55ebb606;
    ram_cell[     693] = 32'h7c1fd646;
    ram_cell[     694] = 32'h6b7e383e;
    ram_cell[     695] = 32'h671bea61;
    ram_cell[     696] = 32'h3ac556c9;
    ram_cell[     697] = 32'h9b73d0e2;
    ram_cell[     698] = 32'hbf54603c;
    ram_cell[     699] = 32'h48736958;
    ram_cell[     700] = 32'hed92041b;
    ram_cell[     701] = 32'haf68f593;
    ram_cell[     702] = 32'h09721286;
    ram_cell[     703] = 32'h1eb087af;
    ram_cell[     704] = 32'h77a891a3;
    ram_cell[     705] = 32'hd0b104be;
    ram_cell[     706] = 32'hc5375778;
    ram_cell[     707] = 32'h71f46ec7;
    ram_cell[     708] = 32'hec5435ac;
    ram_cell[     709] = 32'h6a1017c3;
    ram_cell[     710] = 32'h641e8209;
    ram_cell[     711] = 32'h67ea4cf9;
    ram_cell[     712] = 32'h2f418943;
    ram_cell[     713] = 32'h48b9285f;
    ram_cell[     714] = 32'h2ad03774;
    ram_cell[     715] = 32'hebc08eff;
    ram_cell[     716] = 32'h8d9f79c3;
    ram_cell[     717] = 32'h02613e99;
    ram_cell[     718] = 32'h99f40dc3;
    ram_cell[     719] = 32'h17a7120e;
    ram_cell[     720] = 32'h6d55869c;
    ram_cell[     721] = 32'h8ed7acb5;
    ram_cell[     722] = 32'h3b0f9bef;
    ram_cell[     723] = 32'h12667cf7;
    ram_cell[     724] = 32'h9d4051de;
    ram_cell[     725] = 32'h6227ef03;
    ram_cell[     726] = 32'hb72762a1;
    ram_cell[     727] = 32'hee387558;
    ram_cell[     728] = 32'h614b632e;
    ram_cell[     729] = 32'heebfe446;
    ram_cell[     730] = 32'h8ef758d7;
    ram_cell[     731] = 32'h1a516645;
    ram_cell[     732] = 32'h12d92525;
    ram_cell[     733] = 32'hfb5dd659;
    ram_cell[     734] = 32'h262666dd;
    ram_cell[     735] = 32'h6e35b517;
    ram_cell[     736] = 32'h62d3f583;
    ram_cell[     737] = 32'h6d85407c;
    ram_cell[     738] = 32'h7900f688;
    ram_cell[     739] = 32'heb7b08c3;
    ram_cell[     740] = 32'hbcf145f9;
    ram_cell[     741] = 32'h79b7b9cb;
    ram_cell[     742] = 32'hbc2041e3;
    ram_cell[     743] = 32'h46daba3b;
    ram_cell[     744] = 32'h446676be;
    ram_cell[     745] = 32'h9d7fdac1;
    ram_cell[     746] = 32'h430911f9;
    ram_cell[     747] = 32'ha1e8a918;
    ram_cell[     748] = 32'had08b49f;
    ram_cell[     749] = 32'h881111b7;
    ram_cell[     750] = 32'hc73eea97;
    ram_cell[     751] = 32'hcc17fcf1;
    ram_cell[     752] = 32'hc75763a7;
    ram_cell[     753] = 32'h5d6f4567;
    ram_cell[     754] = 32'h854d7f5e;
    ram_cell[     755] = 32'h59010523;
    ram_cell[     756] = 32'h3478864b;
    ram_cell[     757] = 32'h17fb8f41;
    ram_cell[     758] = 32'h988aca6a;
    ram_cell[     759] = 32'h450ab7c1;
    ram_cell[     760] = 32'h537557f4;
    ram_cell[     761] = 32'hd152efc7;
    ram_cell[     762] = 32'h6c8c6cb6;
    ram_cell[     763] = 32'h447b6b8a;
    ram_cell[     764] = 32'hc3f8fb89;
    ram_cell[     765] = 32'h87457037;
    ram_cell[     766] = 32'h31806b34;
    ram_cell[     767] = 32'ha722afe3;
end

endmodule

